module font_rom ( input [7:0]	addr_ones, addr_tens, addr_hunds, addr_thous,
						output [15:0]	data_ones, data_tens, data_hunds, data_thous
					 );

	parameter ADDR_WIDTH = 8;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:159][15:0] ROM = {
         // code x00
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000011111000000, // 2  *****
        16'b0000110001100000, // 3 **   **
        16'b0000110001100000, // 4 **   **
        16'b0000110011100000, // 5 **  ***
        16'b0000110111100000, // 6 ** ****
        16'b0000111101100000, // 7 **** **
        16'b0000111001100000, // 8 ***  **
        16'b0000110001100000, // 9 **   **
        16'b0000110001100000, // a **   **
        16'b0000011111000000, // b  *****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x01
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000110000000, // 2
        16'b0000001110000000, // 3
        16'b0000011110000000, // 4    **
        16'b0000000110000000, // 5   ***
        16'b0000000110000000, // 6  ****
        16'b0000000110000000, // 7    **
        16'b0000000110000000, // 8    **
        16'b0000000110000000, // 9    **
        16'b0000000110000000, // a    **
        16'b0000011111100000, // b    **
        16'b0000000000000000, // c    **
        16'b0000000000000000, // d  ******
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x02
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000011111000000, // 2  *****
        16'b0000110001100000, // 3 **   **
        16'b0000000001100000, // 4      **
        16'b0000000011000000, // 5     **
        16'b0000000110000000, // 6    **
        16'b0000001100000000, // 7   **
        16'b0000011000000000, // 8  **
        16'b0000110000000000, // 9 **
        16'b0000110001100000, // a **   **
        16'b0000111111100000, // b *******
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x03
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000011111000000, // 2  *****
        16'b0000110001100000, // 3 **   **
        16'b0000000001100000, // 4      **
        16'b0000000001100000, // 5      **
        16'b0000001111000000, // 6   ****
        16'b0000000001100000, // 7      **
        16'b0000000001100000, // 8      **
        16'b0000000001100000, // 9      **
        16'b0000110001100000, // a **   **
        16'b0000011111000000, // b  *****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x04
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000011000000, // 2     **
        16'b0000000111000000, // 3    ***
        16'b0000001111000000, // 4   ****
        16'b0000011011000000, // 5  ** **
        16'b0000110011000000, // 6 **  **
        16'b0000111111100000, // 7 *******
        16'b0000000011000000, // 8     **
        16'b0000000011000000, // 9     **
        16'b0000000011000000, // a     **
        16'b0000000111100000, // b    ****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x05
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000111111100000, // 2 *******
        16'b0000110000000000, // 3 **
        16'b0000110000000000, // 4 **
        16'b0000110000000000, // 5 **
        16'b0000111111000000, // 6 ******
        16'b0000000001100000, // 7      **
        16'b0000000001100000, // 8      **
        16'b0000000001100000, // 9      **
        16'b0000110001100000, // a **   **
        16'b0000011111000000, // b  *****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x06
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000001110000000, // 2   ***
        16'b0000011000000000, // 3  **
        16'b0000110000000000, // 4 **
        16'b0000110000000000, // 5 **
        16'b0000111111000000, // 6 ******
        16'b0000110001100000, // 7 **   **
        16'b0000110001100000, // 8 **   **
        16'b0000110001100000, // 9 **   **
        16'b0000110001100000, // a **   **
        16'b0000011111000000, // b  *****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x07
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000111111100000, // 2 *******
        16'b0000110001100000, // 3 **   **
        16'b0000000001100000, // 4      **
        16'b0000000001100000, // 5      **
        16'b0000000011000000, // 6     **
        16'b0000000110000000, // 7    **
        16'b0000001100000000, // 8   **
        16'b0000001100000000, // 9   **
        16'b0000001100000000, // a   **
        16'b0000001100000000, // b   **
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x08
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000011111000000, // 2  *****
        16'b0000110001100000, // 3 **   **
        16'b0000110001100000, // 4 **   **
        16'b0000110001100000, // 5 **   **
        16'b0000011111000000, // 6  *****
        16'b0000110001100000, // 7 **   **
        16'b0000110001100000, // 8 **   **
        16'b0000110001100000, // 9 **   **
        16'b0000110001100000, // a **   **
        16'b0000011111000000, // b  *****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x09
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000011111000000, // 2  *****
        16'b0000110001100000, // 3 **   **
        16'b0000110001100000, // 4 **   **
        16'b0000110001100000, // 5 **   **
        16'b0000011111100000, // 6  ******
        16'b0000000001100000, // 7      **
        16'b0000000001100000, // 8      **
        16'b0000000001100000, // 9      **
        16'b0000000011000000, // a     **
        16'b0000011110000000, // b  ****
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
        };

	assign data_ones = ROM[addr_ones];
	assign data_tens = ROM[addr_tens];
	assign data_hunds = ROM[addr_hunds];
	assign data_thous = ROM[addr_thous];

endmodule  